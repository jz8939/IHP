** sch_path: /home/Joerdson/IHP-Open-PDK/ihp-sg13g2/libs.tech/xschem/Mixer5GHz.sch
**.subckt Mixer5GHz RFN RFP VDC IFP IFN GND IDC OSCN OSCP VCC ICC GND
*.iopin RFN
*.iopin RFP
*.iopin VDC
*.iopin IFP
*.iopin IFN
*.iopin GND
*.iopin IDC
*.iopin OSCN
*.iopin OSCP
*.iopin VCC
*.iopin ICC
*.iopin GND
XM6 RFN LON net2 GND sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
XRL2 RFN VDC rppd w=4.50e-6 l=3.20e-6 m=1 b=0
XRL1 RFP VDC rppd w=4.50e-6 l=3.20e-6 m=1 b=0
XM8 RFN LOP net3 GND sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
XM7 RFP LON net3 GND sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
XM5 RFP LOP net2 GND sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
XM4 net3 IFN net1 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM3 net2 IFP net1 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM2 IDC IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XM1 net1 IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XM11 LOP LON net4 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM12 LON LOP net4 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM9 IDC IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XM10 net4 IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XC1 VDC LOP cap_cmim w=11.745e-6 l=9.445e-6 m=1
XR1 LOP VDC rppd w=4.4e-6 l=1.5e-6 m=1 b=0
XC2 VDC LON cap_cmim w=11.745e-6 l=9.445e-6 m=1
XR2 LON VDC rppd w=4.4e-6 l=1.5e-6 m=1 b=0
XM13 OSCP OSCN net5 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM14 OSCN OSCP net5 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM15 ICC ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XM16 net5 ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XC3 VCC OSCP cap_cmim w=19.1e-6 l=10.7e-6 m=1
XR3 OSCP VCC rppd w=4.35e-6 l=1.5e-6 m=1 b=0
XC4 VCC OSCN cap_cmim w=19.1e-6 l=10.7e-6 m=1
XR4 OSCN VCC rppd w=4.35e-6 l=1.5e-6 m=1 b=0
L3 VCC OSCP 2.006n m=1
L1 VDC LOP 2.006n m=1
L2 VDC LON 2.006n m=1
L4 VCC OSCN 2.006n m=1
**.ends
.end
