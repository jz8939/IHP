** sch_path: /home/angel/Code/IHP/Mixer5GHz.sch
**.subckt Mixer5GHz RFN RFP VDC IFP IFN GND IDC OSCN OSCP VCC ICC GND
*.iopin RFN
*.iopin RFP
*.iopin VDC
*.iopin IFP
*.iopin IFN
*.iopin GND
*.iopin IDC
*.iopin OSCN
*.iopin OSCP
*.iopin VCC
*.iopin ICC
*.iopin GND
XM6 RFN LON net2 GND sg13_lv_nmos w=60.0u l=0.13u ng=10
XRL2 VDC RFN sub! rppd w=4.50e-6 l=3.20e-6 m=1 b=0
XRL1 VDC RFP sub! rppd w=4.50e-6 l=3.20e-6 m=1 b=0
XM8 RFN LOP net3 GND sg13_lv_nmos w=60.0u l=0.13u ng=10
XM7 RFP LON net3 GND sg13_lv_nmos w=60.0u l=0.13u ng=10
XM5 RFP LOP net2 GND sg13_lv_nmos w=60.0u l=0.13u ng=10
XM4 net3 IFN net1 GND sg13_lv_nmos w=90.0u l=0.13u ng=15
XM3 net2 IFP net1 GND sg13_lv_nmos w=90.0u l=0.13u ng=15
XM2 IDC IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20
XM1 net1 IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20
XM11 LOP LON net4 GND sg13_lv_nmos w=90.0u l=0.13u ng=15
XM12 LON LOP net4 GND sg13_lv_nmos w=90.0u l=0.13u ng=15
XM9 IDC IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20
XM10 net4 IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20
XC1 VDC LOP cap_cmim w=11.745e-6 l=9.445e-6
XR1 VDC LOP sub! rppd w=4.4e-6 l=1.5e-6 m=1 b=0
XC2 VDC LON cap_cmim w=11.745e-6 l=9.445e-6
XR2 VDC LON sub! rppd w=4.4e-6 l=1.5e-6 m=1 b=0
XM13 OSCP OSCN net5 GND sg13_lv_nmos w=90.0u l=0.13u ng=15
XM14 OSCN OSCP net5 GND sg13_lv_nmos w=90.0u l=0.13u ng=15
XM15 ICC ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20
XM16 net5 ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20
XC3 VCC OSCP cap_cmim w=19.1e-6 l=10.7e-6
XR3 VCC OSCP sub! rppd w=4.35e-6 l=1.5e-6 m=1 b=0
XC4 VCC OSCN cap_cmim w=19.1e-6 l=10.7e-6
XR4 VCC OSCN sub! rppd w=4.35e-6 l=1.5e-6 m=1 b=0
L3 VCC OSCP 2.006n
L1 VDC LOP 2.006n
L2 VDC LON 2.006n
L4 VCC OSCN 2.006n
**.ends
.end
